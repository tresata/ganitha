id,x,y
1,1.8858951605446994,0.9604082115601741
2,2.0041264057663586,1.0403196817180977
3,2.166203089543309,0.9216438337721062
4,1.954172979428717,1.1071566582657286
5,2.3314924647036337,0.9677005843374378
6,1.9180772967226227,0.8188749247808329
7,2.0932992502430157,0.8013085715174729
8,1.923195936735381,1.049124293967229
9,1.7383517988067843,0.8994454027942858
10,2.1375166646887163,0.7533985939759434
11,1.9697569304533213,0.9790526216146614
12,1.8628051107434433,0.9528634903011597
13,1.9798743300575612,0.6489056373976361
14,2.4111247138546075,0.6685665540692551
15,2.0822101430371616,0.9663027244053592
16,1.9267805156691795,0.9900682849068371
17,1.8998014184945662,1.3360733744498414
18,1.899215930842022,1.1014630188547376
19,1.9405394796987643,1.1315703415314404
20,1.7861098816704444,1.043370012177357
21,2.0735035815900598,0.9477370259366396
22,1.9913970500652887,1.0216194929544078
23,2.016092377094191,0.9854781282406193
24,2.0395097813887464,1.0874872801645021
25,2.002642389986478,1.0075389114483777
26,1.9321726237377914,1.090383568601841
27,1.8482393903325343,0.8995950441696159
28,1.8593940840087042,0.9650490258105044
29,2.080439151477691,0.9842827120776072
30,2.0566779921292757,0.9768488341726125
31,2.012048353703864,0.9853267684474009
32,1.8326078096645515,0.9187715559918582
33,2.0771151825626304,1.1100610667698592
34,1.719992136334175,1.308657865426066
35,1.954074345758027,0.8709638523654095
36,2.0533607011517976,1.166082035257439
37,2.252556143145334,1.2145586191105706
38,2.1721629981413964,0.7439164121991284
39,2.040112923830971,1.0176434763239897
40,1.9721094742856284,1.0225394604315636
41,1.8065187940659344,0.8144510662116745
42,1.7919207070473129,1.200701280710911
43,2.018839411228971,0.9656926943186231
44,2.085826910216942,1.2401059457556576
45,2.179494467323357,1.155941931546167
46,1.8492210212799765,1.2585994813467494
47,2.1660142600920227,1.1094440060536426
48,2.0508543465581335,1.0608590051558577
49,1.9123740418914328,0.9845613616187958
50,2.0114277772458786,1.0074074967947648
51,0.9759211020360029,1.69284979236148
52,0.9038931728589186,1.1529985992774887
53,0.9857313275561445,1.6615213919892733
54,1.3298422367042948,1.5114546600593544
55,1.0817838520408254,1.5951973403258035
56,1.281552315915003,1.5305330209993808
57,1.1241658686861242,1.2689997872932073
58,0.9804330427555524,1.5395468426615506
59,1.0481669583738003,1.5636478693752003
60,1.1057134596464464,1.4279542595360337
61,1.017685136336627,1.4651387390891666
62,1.1267349832854359,1.7159985324032867
63,0.8269837544461354,1.4427140878805969
64,0.9910531595234036,1.5268198919520335
65,1.2819468971130972,1.608851836555149
66,0.7713255661571558,1.1837952939108851
67,0.8664294473900221,1.6000630598204093
68,1.4875767674243936,1.3638877357352037
69,1.0868757142786842,1.6575638337184977
70,1.0163590182316222,1.1995394407789257
71,0.9202621339009568,1.5461826243833912
72,1.0250611581331974,1.439124019059543
73,0.9829088106458342,1.5191987066907102
74,1.1682126369348178,1.7656159476196938
75,1.1215069258148382,1.734152256733617
76,1.2967305147333177,0.8966366528418429
77,1.3193918131523292,0.94272664092233
78,1.223865051775364,0.9636979929095111
79,1.1443357506155836,0.9494675758691865
80,1.2601135985055956,0.9286271202134427
81,1.2550451485152347,0.6699349491666555
82,1.5558597440207291,0.7530865921814316
83,1.1303154141650262,0.7803672540394107
84,1.2967053554659507,0.9301633586153114
85,1.3221555109341376,0.8272605214991068
86,1.3055897065548119,0.9055519396580074
87,1.3114137975762405,0.9499914729274446
88,1.279749947300198,0.8796302702859775
89,1.2573493152663422,0.8442770992348558
90,1.3203513657409611,0.9696801114545868
91,1.4084067884524023,0.7135641994700725
92,1.3070603965965277,0.7412601794988211
93,1.4299507043689461,0.9130566497914193
94,1.3311062443055866,0.9139265616157835
95,1.30263221221704,1.008917777153598
96,1.2971684824544738,0.9046704392161874
97,1.2960921684394937,0.8747959454301631
98,1.4500170195055047,0.8969129034945627
99,1.2886156529779358,0.9184609824480183
100,1.3047682476996316,0.8687865545989114
101,1.34129162088058,0.9048366196908578
102,1.224932300541484,1.0529202914398095
103,1.2428245395688147,0.8485011603925635
104,1.1507291622389877,0.7886849667728588
105,1.3443334835138283,0.8955119395261486
106,1.2088081898086267,1.1969284841074845
107,1.1506990858536243,1.0066001954922195
108,1.4029319920607721,0.9616450247008271
109,1.2928738426274757,0.9000619010978171
110,1.2167870490819401,1.1231728707426114
111,1.3436778427159757,0.9084873918450035
112,1.3051547752430133,0.8939605841697804
113,1.29392450832213,0.8324116969544083
114,1.3212054713122792,0.9440778967210233
115,1.382979381173592,0.7449325146882393
116,1.3837289287904113,1.0407333880921938
117,1.2268377850362067,0.8974585631313319
118,1.2824414816051848,0.9194196237857746
119,1.2470415229398768,0.8273297928412287
120,1.286020492653493,0.9901271463270676
121,1.3957108932467472,0.6936872858983903
122,1.2308785543192198,0.7828783787643393
123,1.1167065511993455,0.8852329360611296
124,1.3595609348198419,1.0894400711158516
125,1.2703169366257243,0.8543863137404486
126,1.1804280323585112,0.8044959322790964
127,1.4336520121568694,0.9440493423474174
128,1.31480996321265,0.9014314246926426
129,1.0604432164870154,0.8946872292050874
130,1.3263303527900456,0.9091643288257312
131,1.2283407652799254,0.8552557032703055
132,1.3187557756058836,0.8959303207736423
133,1.2827621132872784,0.9442899662870428
134,1.3712193115870845,0.8077148809767868
135,1.197025891759685,0.801636043566108
136,1.2044902788635898,0.8120194537456242
137,1.2117901543802316,0.9469972951087333
138,1.331438723826886,0.896957179124445
139,1.4085777076461814,1.1189006632046448
140,1.5671878633579515,0.9087476549172254
141,1.4043305220298123,0.9410357230796632
142,1.3188488962997067,0.9089748051187261
143,1.2454656119072167,0.9014873504877721
144,1.3996986882144642,1.0243977343975579
145,1.2929193752152381,0.8210186891218625
146,1.4265660562667866,1.0048808104309523
147,1.2692830797706307,0.7189725246442277
148,1.284189803829779,0.9120532958152985
149,1.4255107277050738,0.8535658266873695
150,1.5878378412305891,1.0272252096164451
151,1.9280003118056053,1.660895749545738
152,1.6728886425457836,1.633500198868785
153,1.7925389506719065,1.9803358223662728
154,1.533200995521645,1.9142546231779671
155,1.7500442222897774,1.7317887314385676
156,1.7538080003488146,1.7908585615363948
157,1.7872141234201966,1.4990374442594396
158,1.6598863134730921,1.8744170017518347
159,1.720175475862818,1.5987244599697208
160,1.7689521246922562,1.6917502071570203
161,1.764565937621354,1.7422555749001758
162,1.8541245415377114,1.8012333062734807
163,1.6034147808706356,2.0152885093552793
164,1.7137060107725086,1.745275661717606
165,1.7410714346086695,1.733431667265337
166,1.61211472119022,1.5513351584477224
167,1.6969533160352441,1.8760156869100706
168,1.7609992062564848,1.6535724131012892
169,1.892364499022473,2.190502408118857
170,1.7151986187104933,1.746791136365503
171,1.7559505060698544,1.739045744132873
172,1.8342687148742172,1.5777473280264664
173,1.641410781775027,1.4705329637655336
174,1.7193557262317758,1.7791974087819293
175,1.8763656561032267,1.8029328055283418
176,1.6638511191009175,1.7086147655475057
177,1.7849592461248882,1.7574065602167634
178,1.6231536897328858,1.92228156128578
179,1.6944445619603647,2.1889155267107636
180,1.8871888079977746,1.7652445706087063
181,1.8928418387427928,1.8670809327951778
182,1.6821039306659524,1.742907497679716
183,1.7541601145124135,1.852470536995586
184,1.598537716792164,1.5689957907818328
185,1.9141551679970856,1.6903082045567623
186,1.5646727877629871,1.8825954291703622
187,1.8120949141177782,1.6294050250618621
188,1.716894459608927,1.6602646905150202
189,1.8225866367154429,1.781363645707162
190,1.79250435942207,1.7230789111202187
191,1.732641294040831,1.7581616746235105
192,1.7479554771179617,1.8188540065039973
193,1.8194185970087415,1.5728893841275675
194,1.775482603713787,1.7884952485540617
195,1.8856233241798896,1.756486855880285
196,1.5351746099040917,1.9184730686233002
197,1.751097951642761,1.7657086436568414
198,1.7724479013126908,1.9175295612849328
199,1.695891632234891,1.7340693729487309
200,1.6776703677186495,1.6138847609539213
